class c_180_2;
    rand bit[7:0] data_9_; // rand_mode = ON 

    constraint c1_this    // (constraint_mode = ON) (cb_si.sv:9)
    {
       (data_9_ == 8'hbc);
    }
    constraint c3_this    // (constraint_mode = ON) (cb_si.sv:13)
    {
       (data_9_ != 8'hbc);
    }
endclass

program p_180_2;
    c_180_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz10x1011z1xxz1zx1x1x110xzx11xzzxxzzxxzzxxxzxxxzxzxzzzzzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
