class c_29_2;
    rand bit[7:0] data_8_; // rand_mode = ON 

    constraint c1_this    // (constraint_mode = ON) (cb_si.sv:9)
    {
       (data_8_ == 8'hbc);
    }
    constraint c3_this    // (constraint_mode = ON) (cb_si.sv:13)
    {
       (data_8_ != 8'hbc);
    }
endclass

program p_29_2;
    c_29_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01100z01xzx10z0x00zx10z10xx01011xzzzzzxxzzxxzxxzzxzzzxzxxxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
