class c_83_2;
    rand bit[7:0] data_9_; // rand_mode = ON 

    constraint c1_this    // (constraint_mode = ON) (cb_si.sv:9)
    {
       (data_9_ == 8'hbc);
    }
    constraint c3_this    // (constraint_mode = ON) (cb_si.sv:13)
    {
       (data_9_ != 8'hbc);
    }
endclass

program p_83_2;
    c_83_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00z101zxx0zx10001x00z0xxx101x0xzxzxxzxzxxzxzzxxxzxzzzzzxzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
