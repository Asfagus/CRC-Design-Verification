class cb_scoreboard_illegal extends uvm_scoreboard;
	`uvm_component_utils(cb_scoreboard_illegal)

	uvm_tlm_analysis_fifo #(momsg) message_in_scbd_illegal;

	momsg out;

	function new(string name="cb_scoreboard_illegal",uvm_component parent=null);
		super.new(name, parent);
	endfunction : new

	function void build_phase(uvm_phase phase);
		message_in_scbd_illegal=new("message_in_scbd_illegal",this);
	endfunction: build_phase

	task run_phase(uvm_phase phase);
		fork
			forever begin
				message_in_scbd_illegal.get(out);
				case(out.dataout)
					10'b0010111001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101000110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010101110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101010001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010101101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101010010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010101011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101010100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101000111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010111000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010100111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101011000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010111010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101000101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010110110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101001001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010010111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101101000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010110011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101001100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010011011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101100100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010011101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101100010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010011110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101100001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0010110101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101001010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)

					10'b1001111001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001000110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001101110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001010001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001101101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001010010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001101011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001010100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001000111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001111000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001100111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001011000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001111010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001000101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001110110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001001001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001010111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001101000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001110011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001001100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001011011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001100100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001011101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001100010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001011110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001100001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001110101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001001010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)

					10'b1010111001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010000110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010101110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010010001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010101101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010010010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010101011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010010100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010000111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010111000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010100111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010011000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010111010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010000101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010110110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010001001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010010111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010101000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010110011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010001100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010011011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010100100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010011101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010100010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010011110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010100001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010110101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010001010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)

					10'b1100111001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011000110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100101110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011010001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100101101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011010010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100101011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011010100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011000111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100111000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100100111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011011000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100111010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011000101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100110110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011001001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100010111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011101000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100110011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011001100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100011011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011100100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100011101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011100010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100011110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011100001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100110101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011001010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)

					10'b0100111001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011000110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100101110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011010001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100101101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011010010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100101011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011010100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011000111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100111000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100100111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011011000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100111010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011000101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100110110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011001001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100010111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011101000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100110011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011001100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100011011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011100100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100011101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011100010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100011110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011100001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100110101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011001010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)

					10'b0101111001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101000110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101101110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101010001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101101101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101010010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101101011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101010100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101000111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101111000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101100111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101011000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101111010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101000101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101110110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101001001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101010111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101101000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101110011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101001100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101011011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101100100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101011101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101100010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101011110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101100001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101110101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101001010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)

					10'b0110111001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110000110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110101110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110010001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110101101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110010010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110101011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110010100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110000111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110111000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110100111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110011000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110111010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110000101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110110110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110001001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110010111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110101000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110110011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110001100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110011011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110100100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110011101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110100010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110011110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110100001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110110101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110001010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)

					10'b1000111001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111000110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000101110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111010001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000101101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111010010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000100011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000101011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111010100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000100101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000100110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111000111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000111000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000100111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111011000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000101001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000101010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0001001011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000101100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0001001101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0001001110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000111010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111000101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000110110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111001001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1110110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000110001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1110110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000110010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000010011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1110110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000110100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000010101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000010110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000010111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111101000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000110011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111001100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000011001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000011010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000011011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111100100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000011100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000011101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111100010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000011110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111100001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1000110101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0111001010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					
					10'b0010111100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1101000011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001111100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110000011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010111100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101000011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1100111100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0011000011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0100111100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1011000011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0101111100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1010000011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0110111100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1001000011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0001010111:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1110101000:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0001011011:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1110100100:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0001011101:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1110100010:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b0001011110:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					10'b1110100001:`uvm_info(get_type_name(),$sformatf("legal code act:%h ",out.dataout),UVM_MEDIUM)
					default: `uvm_error("illegal code",$sformatf("Failed act:%h",out.dataout))
				endcase
			end
		join

	endtask: run_phase

endclass: cb_scoreboard_illegal
