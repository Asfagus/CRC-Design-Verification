class c_157_2;
    rand bit[7:0] data_8_; // rand_mode = ON 

    constraint c1_this    // (constraint_mode = ON) (cb_si.sv:9)
    {
       (data_8_ == 8'hbc);
    }
    constraint c3_this    // (constraint_mode = ON) (cb_si.sv:13)
    {
       (data_8_ != 8'hbc);
    }
endclass

program p_157_2;
    c_157_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xzzz0z1x10zxxz010x1x01010x1z01zzxxxzxzzzxzzxxzxxzxzxxxxxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
