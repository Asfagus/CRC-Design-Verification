// This is a message from monout to scorboard1

class momsg;	
	logic startout,pushout;
	logic [9:0] dataout;

endclass:momsg
