// This is a message from monin to scorboard0

class mimsg;	
	logic reset,startin,pushin;
	logic [8:0] datain;

endclass:mimsg
